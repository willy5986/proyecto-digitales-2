module Serial_Paralelo_phy_tx(clk_32f, data_in, default_values, active, idle_out, data_out);